`define ALU_OP_ADD 		5'b00000
`define ALU_OP_SUB 		5'b10000
`define ALU_OP_AND 		5'b00111
`define ALU_OP_OR  		5'b00110
`define ALU_OP_XOR 		5'b00100
`define ALU_OP_MUL 		5'b01000
`define ALU_OP_MULH 	5'b01001
`define ALU_OP_MULHU 	5'b01011
`define ALU_OP_MULHSU 	5'b01010
`define ALU_OP_DIV 		5'b01100
`define ALU_OP_DIVU 	5'b01101
`define ALU_OP_REM 		5'b01110
`define ALU_OP_REMU 	5'b01111
`define ALU_OP_LSH		5'b00001
`define ALU_OP_RSH		5'b00101
`define ALU_OP_ARSH		5'b10101
`define ALU_OP_LESS		5'b00010
`define ALU_OP_LESS_U	5'b00011

`define ALU_OP_PT1		5'b11000
`define ALU_OP_PT2		5'b11001

`define ALU_OPERATION_WIDTH 5
