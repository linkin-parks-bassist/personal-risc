module top();
	instr_decoder instrdec();
endmodule
