`define SRAM_COMMAND_NO_CMD			0
`define SRAM_COMMAND_READ8  		1
`define SRAM_COMMAND_READ16  		3
`define SRAM_COMMAND_READ32  		5
`define SRAM_COMMAND_WRITE8 		2
`define SRAM_COMMAND_WRITE16 		4
`define SRAM_COMMAND_WRITE32 		6

`define SRAM_COMMAND_BITS $clog2(7)
