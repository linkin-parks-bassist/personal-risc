module top();
	
endmodule
